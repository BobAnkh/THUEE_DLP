module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	always @(*)
		case (Address[10:2])
			9'd0:    Instruction <= 32'h08000003;
			9'd1:    Instruction <= 32'h08000172;
			9'd2:    Instruction <= 32'h0800019f;
			9'd3:    Instruction <= 32'h24090014;
			9'd4:    Instruction <= 32'h01200008;
			9'd5:    Instruction <= 32'h0000a021;
			9'd6:    Instruction <= 32'h2008003f;
			9'd7:    Instruction <= 32'hae880000;
			9'd8:    Instruction <= 32'h20080006;
			9'd9:    Instruction <= 32'hae880004;
			9'd10:    Instruction <= 32'h2008005b;
			9'd11:    Instruction <= 32'hae880008;
			9'd12:    Instruction <= 32'h2008004b;
			9'd13:    Instruction <= 32'hae88000c;
			9'd14:    Instruction <= 32'h20080066;
			9'd15:    Instruction <= 32'hae880010;
			9'd16:    Instruction <= 32'h2008006d;
			9'd17:    Instruction <= 32'hae880014;
			9'd18:    Instruction <= 32'h2008007d;
			9'd19:    Instruction <= 32'hae880018;
			9'd20:    Instruction <= 32'h20080007;
			9'd21:    Instruction <= 32'hae88001c;
			9'd22:    Instruction <= 32'h2008007f;
			9'd23:    Instruction <= 32'hae880020;
			9'd24:    Instruction <= 32'h2008006f;
			9'd25:    Instruction <= 32'hae880024;
			9'd26:    Instruction <= 32'h20080077;
			9'd27:    Instruction <= 32'hae880028;
			9'd28:    Instruction <= 32'h2008007c;
			9'd29:    Instruction <= 32'hae88002c;
			9'd30:    Instruction <= 32'h20080039;
			9'd31:    Instruction <= 32'hae880030;
			9'd32:    Instruction <= 32'h2008005e;
			9'd33:    Instruction <= 32'hae880034;
			9'd34:    Instruction <= 32'h20080079;
			9'd35:    Instruction <= 32'hae880038;
			9'd36:    Instruction <= 32'h20080071;
			9'd37:    Instruction <= 32'hae88003c;
			9'd38:    Instruction <= 32'h20083dd6;
			9'd39:    Instruction <= 32'hae880040;
			9'd40:    Instruction <= 32'h20083fc9;
			9'd41:    Instruction <= 32'hae880044;
			9'd42:    Instruction <= 32'h200878c5;
			9'd43:    Instruction <= 32'hae880048;
			9'd44:    Instruction <= 32'h200850c0;
			9'd45:    Instruction <= 32'hae88004c;
			9'd46:    Instruction <= 32'h200818e7;
			9'd47:    Instruction <= 32'hae880050;
			9'd48:    Instruction <= 32'h2008006e;
			9'd49:    Instruction <= 32'hae880054;
			9'd50:    Instruction <= 32'h20085ab4;
			9'd51:    Instruction <= 32'hae880058;
			9'd52:    Instruction <= 32'h200805bb;
			9'd53:    Instruction <= 32'hae88005c;
			9'd54:    Instruction <= 32'h200849a0;
			9'd55:    Instruction <= 32'hae880060;
			9'd56:    Instruction <= 32'h20083282;
			9'd57:    Instruction <= 32'hae880064;
			9'd58:    Instruction <= 32'h200843f1;
			9'd59:    Instruction <= 32'hae880068;
			9'd60:    Instruction <= 32'h20080779;
			9'd61:    Instruction <= 32'hae88006c;
			9'd62:    Instruction <= 32'h200811f4;
			9'd63:    Instruction <= 32'hae880070;
			9'd64:    Instruction <= 32'h20081757;
			9'd65:    Instruction <= 32'hae880074;
			9'd66:    Instruction <= 32'h20086f1a;
			9'd67:    Instruction <= 32'hae880078;
			9'd68:    Instruction <= 32'h2008584b;
			9'd69:    Instruction <= 32'hae88007c;
			9'd70:    Instruction <= 32'h20084fd2;
			9'd71:    Instruction <= 32'hae880080;
			9'd72:    Instruction <= 32'h20083989;
			9'd73:    Instruction <= 32'hae880084;
			9'd74:    Instruction <= 32'h200873a5;
			9'd75:    Instruction <= 32'hae880088;
			9'd76:    Instruction <= 32'h20084d19;
			9'd77:    Instruction <= 32'hae88008c;
			9'd78:    Instruction <= 32'h2008015d;
			9'd79:    Instruction <= 32'hae880090;
			9'd80:    Instruction <= 32'h20082ab6;
			9'd81:    Instruction <= 32'hae880094;
			9'd82:    Instruction <= 32'h20084b83;
			9'd83:    Instruction <= 32'hae880098;
			9'd84:    Instruction <= 32'h200802f7;
			9'd85:    Instruction <= 32'hae88009c;
			9'd86:    Instruction <= 32'h20083f59;
			9'd87:    Instruction <= 32'hae8800a0;
			9'd88:    Instruction <= 32'h20085adb;
			9'd89:    Instruction <= 32'hae8800a4;
			9'd90:    Instruction <= 32'h20081093;
			9'd91:    Instruction <= 32'hae8800a8;
			9'd92:    Instruction <= 32'h2008547c;
			9'd93:    Instruction <= 32'hae8800ac;
			9'd94:    Instruction <= 32'h20085925;
			9'd95:    Instruction <= 32'hae8800b0;
			9'd96:    Instruction <= 32'h20081a25;
			9'd97:    Instruction <= 32'hae8800b4;
			9'd98:    Instruction <= 32'h20083c3b;
			9'd99:    Instruction <= 32'hae8800b8;
			9'd100:    Instruction <= 32'h200875ed;
			9'd101:    Instruction <= 32'hae8800bc;
			9'd102:    Instruction <= 32'h20087fd3;
			9'd103:    Instruction <= 32'hae8800c0;
			9'd104:    Instruction <= 32'h2008604e;
			9'd105:    Instruction <= 32'hae8800c4;
			9'd106:    Instruction <= 32'h20087d0c;
			9'd107:    Instruction <= 32'hae8800c8;
			9'd108:    Instruction <= 32'h200808aa;
			9'd109:    Instruction <= 32'hae8800cc;
			9'd110:    Instruction <= 32'h20085802;
			9'd111:    Instruction <= 32'hae8800d0;
			9'd112:    Instruction <= 32'h20087e4a;
			9'd113:    Instruction <= 32'hae8800d4;
			9'd114:    Instruction <= 32'h20086b2f;
			9'd115:    Instruction <= 32'hae8800d8;
			9'd116:    Instruction <= 32'h20084dd1;
			9'd117:    Instruction <= 32'hae8800dc;
			9'd118:    Instruction <= 32'h20084b83;
			9'd119:    Instruction <= 32'hae8800e0;
			9'd120:    Instruction <= 32'h200807ef;
			9'd121:    Instruction <= 32'hae8800e4;
			9'd122:    Instruction <= 32'h20085d0f;
			9'd123:    Instruction <= 32'hae8800e8;
			9'd124:    Instruction <= 32'h20086b21;
			9'd125:    Instruction <= 32'hae8800ec;
			9'd126:    Instruction <= 32'h20085896;
			9'd127:    Instruction <= 32'hae8800f0;
			9'd128:    Instruction <= 32'h200878b6;
			9'd129:    Instruction <= 32'hae8800f4;
			9'd130:    Instruction <= 32'h20081db8;
			9'd131:    Instruction <= 32'hae8800f8;
			9'd132:    Instruction <= 32'h20086330;
			9'd133:    Instruction <= 32'hae8800fc;
			9'd134:    Instruction <= 32'h200840bf;
			9'd135:    Instruction <= 32'hae880100;
			9'd136:    Instruction <= 32'h20081e14;
			9'd137:    Instruction <= 32'hae880104;
			9'd138:    Instruction <= 32'h20084368;
			9'd139:    Instruction <= 32'hae880108;
			9'd140:    Instruction <= 32'h20081e5a;
			9'd141:    Instruction <= 32'hae88010c;
			9'd142:    Instruction <= 32'h200805f6;
			9'd143:    Instruction <= 32'hae880110;
			9'd144:    Instruction <= 32'h20085977;
			9'd145:    Instruction <= 32'hae880114;
			9'd146:    Instruction <= 32'h20080e13;
			9'd147:    Instruction <= 32'hae880118;
			9'd148:    Instruction <= 32'h20087d25;
			9'd149:    Instruction <= 32'hae88011c;
			9'd150:    Instruction <= 32'h20084d8e;
			9'd151:    Instruction <= 32'hae880120;
			9'd152:    Instruction <= 32'h2008418d;
			9'd153:    Instruction <= 32'hae880124;
			9'd154:    Instruction <= 32'h20087384;
			9'd155:    Instruction <= 32'hae880128;
			9'd156:    Instruction <= 32'h200870b8;
			9'd157:    Instruction <= 32'hae88012c;
			9'd158:    Instruction <= 32'h200816c6;
			9'd159:    Instruction <= 32'hae880130;
			9'd160:    Instruction <= 32'h20087fc1;
			9'd161:    Instruction <= 32'hae880134;
			9'd162:    Instruction <= 32'h20086848;
			9'd163:    Instruction <= 32'hae880138;
			9'd164:    Instruction <= 32'h200805c2;
			9'd165:    Instruction <= 32'hae88013c;
			9'd166:    Instruction <= 32'h200872cf;
			9'd167:    Instruction <= 32'hae880140;
			9'd168:    Instruction <= 32'h2008200a;
			9'd169:    Instruction <= 32'hae880144;
			9'd170:    Instruction <= 32'h20084740;
			9'd171:    Instruction <= 32'hae880148;
			9'd172:    Instruction <= 32'h20081fad;
			9'd173:    Instruction <= 32'hae88014c;
			9'd174:    Instruction <= 32'h20080e83;
			9'd175:    Instruction <= 32'hae880150;
			9'd176:    Instruction <= 32'h20084261;
			9'd177:    Instruction <= 32'hae880154;
			9'd178:    Instruction <= 32'h2008366c;
			9'd179:    Instruction <= 32'hae880158;
			9'd180:    Instruction <= 32'h20086643;
			9'd181:    Instruction <= 32'hae88015c;
			9'd182:    Instruction <= 32'h2008127f;
			9'd183:    Instruction <= 32'hae880160;
			9'd184:    Instruction <= 32'h200831f4;
			9'd185:    Instruction <= 32'hae880164;
			9'd186:    Instruction <= 32'h2008582d;
			9'd187:    Instruction <= 32'hae880168;
			9'd188:    Instruction <= 32'h20086ffd;
			9'd189:    Instruction <= 32'hae88016c;
			9'd190:    Instruction <= 32'h20085687;
			9'd191:    Instruction <= 32'hae880170;
			9'd192:    Instruction <= 32'h20081b5f;
			9'd193:    Instruction <= 32'hae880174;
			9'd194:    Instruction <= 32'h20085abb;
			9'd195:    Instruction <= 32'hae880178;
			9'd196:    Instruction <= 32'h20087553;
			9'd197:    Instruction <= 32'hae88017c;
			9'd198:    Instruction <= 32'h20086861;
			9'd199:    Instruction <= 32'hae880180;
			9'd200:    Instruction <= 32'h20086e1d;
			9'd201:    Instruction <= 32'hae880184;
			9'd202:    Instruction <= 32'h200835bd;
			9'd203:    Instruction <= 32'hae880188;
			9'd204:    Instruction <= 32'h20087bbc;
			9'd205:    Instruction <= 32'hae88018c;
			9'd206:    Instruction <= 32'h20085d62;
			9'd207:    Instruction <= 32'hae880190;
			9'd208:    Instruction <= 32'h20087580;
			9'd209:    Instruction <= 32'hae880194;
			9'd210:    Instruction <= 32'h20085250;
			9'd211:    Instruction <= 32'hae880198;
			9'd212:    Instruction <= 32'h200811c1;
			9'd213:    Instruction <= 32'hae88019c;
			9'd214:    Instruction <= 32'h20083865;
			9'd215:    Instruction <= 32'hae8801a0;
			9'd216:    Instruction <= 32'h200864fa;
			9'd217:    Instruction <= 32'hae8801a4;
			9'd218:    Instruction <= 32'h20081dab;
			9'd219:    Instruction <= 32'hae8801a8;
			9'd220:    Instruction <= 32'h20087945;
			9'd221:    Instruction <= 32'hae8801ac;
			9'd222:    Instruction <= 32'h20085620;
			9'd223:    Instruction <= 32'hae8801b0;
			9'd224:    Instruction <= 32'h20081c08;
			9'd225:    Instruction <= 32'hae8801b4;
			9'd226:    Instruction <= 32'h200831cd;
			9'd227:    Instruction <= 32'hae8801b8;
			9'd228:    Instruction <= 32'h200814b8;
			9'd229:    Instruction <= 32'hae8801bc;
			9'd230:    Instruction <= 32'h20085d99;
			9'd231:    Instruction <= 32'hae8801c0;
			9'd232:    Instruction <= 32'h20086c9d;
			9'd233:    Instruction <= 32'hae8801c4;
			9'd234:    Instruction <= 32'h200827aa;
			9'd235:    Instruction <= 32'hae8801c8;
			9'd236:    Instruction <= 32'h200872a1;
			9'd237:    Instruction <= 32'hae8801cc;
			9'd238:    Instruction <= 32'h2008533f;
			9'd239:    Instruction <= 32'hae8801d0;
			9'd240:    Instruction <= 32'h20086cc2;
			9'd241:    Instruction <= 32'hae8801d4;
			9'd242:    Instruction <= 32'h20080e41;
			9'd243:    Instruction <= 32'hae8801d8;
			9'd244:    Instruction <= 32'h20086c6a;
			9'd245:    Instruction <= 32'hae8801dc;
			9'd246:    Instruction <= 32'h20082981;
			9'd247:    Instruction <= 32'hae8801e0;
			9'd248:    Instruction <= 32'h20085783;
			9'd249:    Instruction <= 32'hae8801e4;
			9'd250:    Instruction <= 32'h2008748d;
			9'd251:    Instruction <= 32'hae8801e8;
			9'd252:    Instruction <= 32'h20083e81;
			9'd253:    Instruction <= 32'hae8801ec;
			9'd254:    Instruction <= 32'h20085c13;
			9'd255:    Instruction <= 32'hae8801f0;
			9'd256:    Instruction <= 32'h2008478e;
			9'd257:    Instruction <= 32'hae8801f4;
			9'd258:    Instruction <= 32'h200867f4;
			9'd259:    Instruction <= 32'hae8801f8;
			9'd260:    Instruction <= 32'h20086bf4;
			9'd261:    Instruction <= 32'hae8801fc;
			9'd262:    Instruction <= 32'h20082c17;
			9'd263:    Instruction <= 32'hae880200;
			9'd264:    Instruction <= 32'h20082126;
			9'd265:    Instruction <= 32'hae880204;
			9'd266:    Instruction <= 32'h20085004;
			9'd267:    Instruction <= 32'hae880208;
			9'd268:    Instruction <= 32'h20087fa6;
			9'd269:    Instruction <= 32'hae88020c;
			9'd270:    Instruction <= 32'h20083d2a;
			9'd271:    Instruction <= 32'hae880210;
			9'd272:    Instruction <= 32'h2008143f;
			9'd273:    Instruction <= 32'hae880214;
			9'd274:    Instruction <= 32'h20082b3e;
			9'd275:    Instruction <= 32'hae880218;
			9'd276:    Instruction <= 32'h20084a73;
			9'd277:    Instruction <= 32'hae88021c;
			9'd278:    Instruction <= 32'h20087ef4;
			9'd279:    Instruction <= 32'hae880220;
			9'd280:    Instruction <= 32'h2008141f;
			9'd281:    Instruction <= 32'hae880224;
			9'd282:    Instruction <= 32'h200850a3;
			9'd283:    Instruction <= 32'hae880228;
			9'd284:    Instruction <= 32'h200875a4;
			9'd285:    Instruction <= 32'hae88022c;
			9'd286:    Instruction <= 32'h20083a25;
			9'd287:    Instruction <= 32'hae880230;
			9'd288:    Instruction <= 32'h20080f93;
			9'd289:    Instruction <= 32'hae880234;
			9'd290:    Instruction <= 32'h2008591d;
			9'd291:    Instruction <= 32'hae880238;
			9'd292:    Instruction <= 32'h20082578;
			9'd293:    Instruction <= 32'hae88023c;
			9'd294:    Instruction <= 32'h3c014000;
			9'd295:    Instruction <= 32'h34340008;
			9'd296:    Instruction <= 32'h20080000;
			9'd297:    Instruction <= 32'hae880000;
			9'd298:    Instruction <= 32'h2295fffc;
			9'd299:    Instruction <= 32'h2008ff9b;
			9'd300:    Instruction <= 32'haea80000;
			9'd301:    Instruction <= 32'h2295fff8;
			9'd302:    Instruction <= 32'h2008ff9b;
			9'd303:    Instruction <= 32'haea80000;
			9'd304:    Instruction <= 32'h201d0400;
			9'd305:    Instruction <= 32'h3c014000;
			9'd306:    Instruction <= 32'h34350014;
			9'd307:    Instruction <= 32'h8eb60000;
			9'd308:    Instruction <= 32'h24100040;
			9'd309:    Instruction <= 32'h24110080;
			9'd310:    Instruction <= 32'h00102021;
			9'd311:    Instruction <= 32'h00112821;
			9'd312:    Instruction <= 32'h0c000150;
			9'd313:    Instruction <= 32'h8ea80000;
			9'd314:    Instruction <= 32'h01161022;
			9'd315:    Instruction <= 32'h20090080;
			9'd316:    Instruction <= 32'h200a0040;
			9'd317:    Instruction <= 32'h11200004;
			9'd318:    Instruction <= 32'h2129ffff;
			9'd319:    Instruction <= 32'h8d4b0000;
			9'd320:    Instruction <= 32'h214a0004;
			9'd321:    Instruction <= 32'h0800013d;
			9'd322:    Instruction <= 32'h20080003;
			9'd323:    Instruction <= 32'hae880000;
			9'd324:    Instruction <= 32'h3c014000;
			9'd325:    Instruction <= 32'h34350010;
			9'd326:    Instruction <= 32'h20160000;
			9'd327:    Instruction <= 32'h1000ffff;
			9'd328:    Instruction <= 32'h00054080;
			9'd329:    Instruction <= 32'h01044020;
			9'd330:    Instruction <= 32'h8d090000;
			9'd331:    Instruction <= 32'h8d0a0004;
			9'd332:    Instruction <= 32'had0a0000;
			9'd333:    Instruction <= 32'had090004;
			9'd334:    Instruction <= 32'h00001021;
			9'd335:    Instruction <= 32'h03e00008;
			9'd336:    Instruction <= 32'h23bdfff4;
			9'd337:    Instruction <= 32'hafbf0000;
			9'd338:    Instruction <= 32'hafb00004;
			9'd339:    Instruction <= 32'hafb10008;
			9'd340:    Instruction <= 32'h00049021;
			9'd341:    Instruction <= 32'h00059821;
			9'd342:    Instruction <= 32'h24100000;
			9'd343:    Instruction <= 32'h0213402a;
			9'd344:    Instruction <= 32'h11000013;
			9'd345:    Instruction <= 32'h2211ffff;
			9'd346:    Instruction <= 32'h0220482a;
			9'd347:    Instruction <= 32'h34010001;
			9'd348:    Instruction <= 32'h00294823;
			9'd349:    Instruction <= 32'h1120000c;
			9'd350:    Instruction <= 32'h00115080;
			9'd351:    Instruction <= 32'h024a5020;
			9'd352:    Instruction <= 32'h8d4b0000;
			9'd353:    Instruction <= 32'h8d4c0004;
			9'd354:    Instruction <= 32'h018b502a;
			9'd355:    Instruction <= 32'h012a4824;
			9'd356:    Instruction <= 32'h11200005;
			9'd357:    Instruction <= 32'h00122021;
			9'd358:    Instruction <= 32'h00112821;
			9'd359:    Instruction <= 32'h0c000148;
			9'd360:    Instruction <= 32'h2231ffff;
			9'd361:    Instruction <= 32'h0800015a;
			9'd362:    Instruction <= 32'h22100001;
			9'd363:    Instruction <= 32'h08000157;
			9'd364:    Instruction <= 32'h8fb10008;
			9'd365:    Instruction <= 32'h8fb00004;
			9'd366:    Instruction <= 32'h8fbf0000;
			9'd367:    Instruction <= 32'h23bd000c;
			9'd368:    Instruction <= 32'h00001021;
			9'd369:    Instruction <= 32'h03e00008;
			9'd370:    Instruction <= 32'h200d0001;
			9'd371:    Instruction <= 32'hae8d0000;
			9'd372:    Instruction <= 32'h2419000f;
			9'd373:    Instruction <= 32'h0002b821;
			9'd374:    Instruction <= 32'h02f96824;
			9'd375:    Instruction <= 32'h0017b902;
			9'd376:    Instruction <= 32'h02f97024;
			9'd377:    Instruction <= 32'h0017b902;
			9'd378:    Instruction <= 32'h02f97824;
			9'd379:    Instruction <= 32'h0017b902;
			9'd380:    Instruction <= 32'h02f9c024;
			9'd381:    Instruction <= 32'h20170000;
			9'd382:    Instruction <= 32'h02d9b024;
			9'd383:    Instruction <= 32'h12c00006;
			9'd384:    Instruction <= 32'h20190004;
			9'd385:    Instruction <= 32'h12d90009;
			9'd386:    Instruction <= 32'h20190008;
			9'd387:    Instruction <= 32'h12d9000c;
			9'd388:    Instruction <= 32'h2019000c;
			9'd389:    Instruction <= 32'h12d9000f;
			9'd390:    Instruction <= 32'h000d6880;
			9'd391:    Instruction <= 32'h01b76820;
			9'd392:    Instruction <= 32'h8db90000;
			9'd393:    Instruction <= 32'h23390800;
			9'd394:    Instruction <= 32'h0800019a;
			9'd395:    Instruction <= 32'h000e7080;
			9'd396:    Instruction <= 32'h01d77020;
			9'd397:    Instruction <= 32'h8dd90000;
			9'd398:    Instruction <= 32'h23390400;
			9'd399:    Instruction <= 32'h0800019a;
			9'd400:    Instruction <= 32'h000f7880;
			9'd401:    Instruction <= 32'h01f77820;
			9'd402:    Instruction <= 32'h8df90000;
			9'd403:    Instruction <= 32'h23390200;
			9'd404:    Instruction <= 32'h0800019a;
			9'd405:    Instruction <= 32'h0018c080;
			9'd406:    Instruction <= 32'h0317c020;
			9'd407:    Instruction <= 32'h8f190000;
			9'd408:    Instruction <= 32'h23390100;
			9'd409:    Instruction <= 32'h0800019a;
			9'd410:    Instruction <= 32'haeb90000;
			9'd411:    Instruction <= 32'h22d60004;
			9'd412:    Instruction <= 32'h20190003;
			9'd413:    Instruction <= 32'hae990000;
			9'd414:    Instruction <= 32'h03400008;
			9'd415:    Instruction <= 32'h1000ffff;
			default:  Instruction <= 32'h0;
		endcase
		
endmodule
